library verilog;
use verilog.vl_types.all;
entity \muddlib07__flopr_c_1x\ is
    port(
        ph1             : in     vl_logic;
        ph2             : in     vl_logic;
        d               : in     vl_logic;
        resetb          : in     vl_logic;
        q               : out    vl_logic;
        vdd             : in     vl_logic;
        gnd             : in     vl_logic
    );
end \muddlib07__flopr_c_1x\;
