library verilog;
use verilog.vl_types.all;
entity \wordlib8__adder_8\ is
    port(
        a               : in     vl_logic_vector(7 downto 0);
        b               : in     vl_logic_vector(7 downto 0);
        cin             : in     vl_logic;
        cout            : out    vl_logic;
        s               : out    vl_logic_vector(7 downto 0);
        vdd             : in     vl_logic;
        vdd_1           : in     vl_logic;
        vdd_1_1         : in     vl_logic;
        vdd_2           : in     vl_logic;
        vdd_3           : in     vl_logic;
        vdd_4           : in     vl_logic;
        vdd_5           : in     vl_logic;
        vdd_6           : in     vl_logic;
        gnd             : in     vl_logic;
        gnd_1           : in     vl_logic;
        gnd_1_1         : in     vl_logic;
        gnd_2           : in     vl_logic;
        gnd_3           : in     vl_logic;
        gnd_4           : in     vl_logic;
        gnd_5           : in     vl_logic;
        gnd_6           : in     vl_logic
    );
end \wordlib8__adder_8\;
