library verilog;
use verilog.vl_types.all;
entity \muddlib07__invbuf_4x\ is
    port(
        s               : in     vl_logic;
        s_out           : out    vl_logic;
        sb_out          : out    vl_logic;
        vdd             : in     vl_logic;
        gnd             : in     vl_logic
    );
end \muddlib07__invbuf_4x\;
