library verilog;
use verilog.vl_types.all;
entity \muddlib07__clkinvbufdual_4x\ is
    port(
        ph1             : in     vl_logic;
        ph2             : in     vl_logic;
        ph1b            : out    vl_logic;
        ph1buf          : out    vl_logic;
        ph2b            : out    vl_logic;
        ph2buf          : out    vl_logic;
        vdd             : in     vl_logic;
        gnd             : in     vl_logic
    );
end \muddlib07__clkinvbufdual_4x\;
