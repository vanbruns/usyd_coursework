library verilog;
use verilog.vl_types.all;
entity \muddlib07__mux2_c_1x\ is
    port(
        d0              : in     vl_logic;
        d1              : in     vl_logic;
        s               : in     vl_logic;
        y               : out    vl_logic;
        vdd             : in     vl_logic;
        gnd             : in     vl_logic
    );
end \muddlib07__mux2_c_1x\;
