library verilog;
use verilog.vl_types.all;
entity \muddpads13_ami05__pad_out\ is
    port(
        dout            : in     vl_logic;
        pad             : out    vl_logic;
        vdd             : in     vl_logic;
        gnd             : in     vl_logic
    );
end \muddpads13_ami05__pad_out\;
