library verilog;
use verilog.vl_types.all;
entity \muddpads13_ami05__pad_corner\ is
    port(
        vdd             : in     vl_logic;
        gnd             : in     vl_logic
    );
end \muddpads13_ami05__pad_corner\;
