library verilog;
use verilog.vl_types.all;
entity \muddpads13_ami05__pad_raw\ is
    port(
        pad             : in     vl_logic;
        vdd             : in     vl_logic;
        gnd             : in     vl_logic
    );
end \muddpads13_ami05__pad_raw\;
