library verilog;
use verilog.vl_types.all;
entity \mips8_vb__regram0\ is
    port(
        read1           : in     vl_logic;
        read2           : in     vl_logic;
        r1              : out    vl_logic;
        r2              : out    vl_logic;
        gnd             : in     vl_logic
    );
end \mips8_vb__regram0\;
