library verilog;
use verilog.vl_types.all;
entity \muddlib07__clkinvbuf_4x\ is
    port(
        ph              : out    vl_logic;
        phb             : out    vl_logic;
        phbuf           : out    vl_logic;
        vdd             : in     vl_logic;
        gnd             : in     vl_logic
    );
end \muddlib07__clkinvbuf_4x\;
