library verilog;
use verilog.vl_types.all;
entity mips_vb_sv_unit is
end mips_vb_sv_unit;
