library verilog;
use verilog.vl_types.all;
entity \muddlib07__mux4_dp_1x\ is
    port(
        d0              : in     vl_logic;
        d1              : in     vl_logic;
        d2              : in     vl_logic;
        d3              : in     vl_logic;
        s0              : in     vl_logic;
        s0b             : in     vl_logic;
        s1              : in     vl_logic;
        s1b             : in     vl_logic;
        y               : out    vl_logic;
        vdd             : in     vl_logic;
        gnd             : in     vl_logic
    );
end \muddlib07__mux4_dp_1x\;
